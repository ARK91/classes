module testbench();


endmodule
