`timescale 1ns/1ns

interface memory_interface(...);


endinterface
