module intro();

   initial $display("======Welcome to UC Santa Cruz Extension======");

   initial begin
      //Display your message here
      $display("Welcome to Verilog");
   end
endmodule
