interface switch_interface(input clk);

    logic [47:0] src_addr;
    logic [31:0] src_data;

endinterface
