interface counter_interface(...);

  // <insert code here>

endinterface

