// File: 4bit_adder_tb.v
// John Hubbard, 23 Jan 2015
// hw1 assignment for UCSC 30207: Digital Design with FPGA

`timescale 1ns/1ns

module add4_tb();
    reg [3:0]a;
    reg [3:0]b;
    wire [4:0]sum;

    add4(a, b, sum);

    initial
    begin
        for (

    end
endmodule

