module packet();
  class packet;
  // <insert you code here>
  endclass
endmodule
