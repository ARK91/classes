// File: 4bit_adder.v
// John Hubbard, 23 Jan 2015
// hw1 assignment for UCSC 30207: Digital Design with FPGA

module add4(a, b, sum);
    input a, b;
    output sum;

    wire [3:0]a;
    wire [3:0]b;
    wire [4:0]sum;

    assign sum = a + b;
endmodule

module add4_struct(a, b, sum);
    input a, b;
    output sum;

    wire [3:0]a;
    wire [3:0]b;
    wire [4:0]sum;

    assign sum[0] = (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]);


    assign sum[1] = (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) +
    (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) +
    (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) +
    (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) +
    (a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]);


    assign sum[2] = (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) +
    (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) +
    (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) +
    (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) +
    (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) +
    (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]);


    assign sum[3] = (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) +
    (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) +
    (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) +
    (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) +
    (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) +
    (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) +
    (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]);


    assign sum[4] =
    (!a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (!a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (!a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&!a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&!a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&!a[0]) & (b[3]&b[2]&b[1]&b[0]) +
    (a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (!b[3]&b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&!b[2]&b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&!b[1]&b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&!b[0]) + (a[3]&a[2]&a[1]&a[0]) & (b[3]&b[2]&b[1]&b[0]);

endmodule
