`timescale 1ns/1ns

program testcase();

endprogram
