class packet;
    rand bit [47:0] src_addr;
    rand bit [31:0] src_data;

    function new();

    endfunction

endclass
