module testbench();



endmodule
