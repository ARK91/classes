module testbench;

  wire        clk;

// Instantiate interface here 

// Instantiate memory design here

// Instantiate testcase here

endmodule
